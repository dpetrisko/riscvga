@00000000
93 00 50 00 13 01 F0 FF 93 01 90 00 13 02 C0 09 
93 02 30 FD 13 03 B0 07 93 03 40 00 33 84 20 00 
B3 84 51 00 33 05 62 00 B3 A5 20 00 33 26 11 00 
B3 36 11 00 33 B7 20 00 B3 77 62 00 33 68 62 00 
B3 C8 22 00 33 99 11 00 B3 D9 72 00 33 0A 62 40 
B3 DA 22 40 6F 00 00 00 13 00 00 00 
