`define IMEM_DEBUG 1
`define DMEM_DEBUG 1
`define INST_DEBUG 1
