@00000000
37 05 00 00 13 05 05 00 37 06 00 10 83 05 05 00 
63 8C 05 00 23 20 B6 00 13 05 15 00 6F F0 1F FF 
6D 79 74 65 73 74 00 00 93 05 E0 02 23 20 B6 00 
23 20 B6 00 B7 80 FF FF 13 01 00 00 B3 D1 20 00 
B7 8E FF FF 13 0E 20 00 63 94 D1 5B B7 80 FF FF 
13 01 10 00 B3 D1 20 00 B7 CE FF 7F 13 0E 30 00 
63 98 D1 59 B7 80 FF FF 13 01 70 00 B3 D1 20 00 
B7 0E 00 02 93 8E 0E F0 13 0E 40 00 63 9A D1 57 
B7 80 FF FF 13 01 E0 00 B3 D1 20 00 B7 0E 04 00 
93 8E EE FF 13 0E 50 00 63 9C D1 55 B7 80 FF FF 
93 80 10 00 13 01 F0 00 B3 D1 20 00 B7 0E 02 00 
93 8E FE FF 13 0E 60 00 63 9C D1 53 93 00 F0 FF 
13 01 00 00 B3 D1 20 00 93 0E F0 FF 13 0E 70 00 
63 90 D1 53 93 00 F0 FF 13 01 10 00 B3 D1 20 00 
B7 0E 00 80 93 8E FE FF 13 0E 80 00 63 92 D1 51 
93 00 F0 FF 13 01 70 00 B3 D1 20 00 B7 0E 00 02 
93 8E FE FF 13 0E 90 00 63 94 D1 4F 93 00 F0 FF 
13 01 E0 00 B3 D1 20 00 B7 0E 04 00 93 8E FE FF 
13 0E A0 00 63 96 D1 4D 93 00 F0 FF 13 01 F0 01 
B3 D1 20 00 93 0E 10 00 13 0E B0 00 63 9A D1 4B 
B7 20 21 21 93 80 10 12 13 01 00 00 B3 D1 20 00 
B7 2E 21 21 93 8E 1E 12 13 0E C0 00 63 9A D1 49 
B7 20 21 21 93 80 10 12 13 01 10 00 B3 D1 20 00 
B7 9E 90 10 93 8E 0E 09 13 0E D0 00 63 9A D1 47 
B7 20 21 21 93 80 10 12 13 01 70 00 B3 D1 20 00 
B7 4E 42 00 93 8E 2E 24 13 0E E0 00 63 9A D1 45 
B7 20 21 21 93 80 10 12 13 01 E0 00 B3 D1 20 00 
B7 8E 00 00 93 8E 4E 48 13 0E F0 00 63 9A D1 43 
B7 20 21 21 93 80 10 12 13 01 F0 01 B3 D1 20 00 
93 0E 00 00 13 0E 00 01 63 9C D1 41 B7 20 21 21 
93 80 10 12 13 01 00 FE B3 D1 20 00 B7 2E 21 21 
93 8E 1E 12 13 0E 10 01 63 9C D1 3F B7 20 21 21 
93 80 10 12 13 01 10 FE B3 D1 20 00 B7 9E 90 10 
93 8E 0E 09 13 0E 20 01 63 9C D1 3D B7 20 21 21 
93 80 10 12 13 01 70 FE B3 D1 20 00 B7 4E 42 00 
93 8E 2E 24 13 0E 30 01 63 9C D1 3B B7 20 21 21 
93 80 10 12 13 01 E0 FE B3 D1 20 00 B7 8E 00 00 
93 8E 4E 48 13 0E 40 01 63 9C D1 39 B7 20 21 21 
93 80 10 12 13 01 F0 FF B3 D1 20 00 93 0E 00 00 
13 0E 50 01 63 9E D1 37 B7 80 FF FF 13 01 10 00 
B3 D0 20 00 B7 CE FF 7F 13 0E 60 01 63 92 D0 37 
B7 80 FF FF 13 01 E0 00 33 D1 20 00 B7 0E 04 00 
93 8E EE FF 13 0E 70 01 63 14 D1 35 93 00 70 00 
B3 D0 10 00 93 0E 00 00 13 0E 80 01 63 9A D0 33 
13 02 00 00 B7 80 FF FF 13 01 10 00 B3 D1 20 00 
13 83 01 00 13 02 12 00 93 02 20 00 E3 14 52 FE 
B7 CE FF 7F 13 0E 90 01 63 14 D3 31 13 02 00 00 
B7 80 FF FF 13 01 E0 00 B3 D1 20 00 13 00 00 00 
13 83 01 00 13 02 12 00 93 02 20 00 E3 12 52 FE 
B7 0E 04 00 93 8E EE FF 13 0E A0 01 63 1A D3 2D 
13 02 00 00 B7 80 FF FF 13 01 F0 00 B3 D1 20 00 
13 00 00 00 13 00 00 00 13 83 01 00 13 02 12 00 
93 02 20 00 E3 10 52 FE B7 0E 02 00 93 8E FE FF 
13 0E B0 01 63 1E D3 29 13 02 00 00 B7 80 FF FF 
13 01 10 00 B3 D1 20 00 13 02 12 00 93 02 20 00 
E3 16 52 FE B7 CE FF 7F 13 0E C0 01 63 9A D1 27 
13 02 00 00 B7 80 FF FF 13 01 70 00 13 00 00 00 
B3 D1 20 00 13 02 12 00 93 02 20 00 E3 14 52 FE 
B7 0E 00 02 93 8E 0E F0 13 0E D0 01 63 92 D1 25 
13 02 00 00 B7 80 FF FF 13 01 F0 00 13 00 00 00 
13 00 00 00 B3 D1 20 00 13 02 12 00 93 02 20 00 
E3 12 52 FE B7 0E 02 00 93 8E FE FF 13 0E E0 01 
63 98 D1 21 13 02 00 00 B7 80 FF FF 13 00 00 00 
13 01 10 00 B3 D1 20 00 13 02 12 00 93 02 20 00 
E3 14 52 FE B7 CE FF 7F 13 0E F0 01 63 92 D1 1F 
13 02 00 00 B7 80 FF FF 13 00 00 00 13 01 70 00 
13 00 00 00 B3 D1 20 00 13 02 12 00 93 02 20 00 
E3 12 52 FE B7 0E 00 02 93 8E 0E F0 13 0E 00 02 
63 98 D1 1B 13 02 00 00 B7 80 FF FF 13 00 00 00 
13 00 00 00 13 01 F0 00 B3 D1 20 00 13 02 12 00 
93 02 20 00 E3 12 52 FE B7 0E 02 00 93 8E FE FF 
13 0E 10 02 63 9E D1 17 13 02 00 00 13 01 10 00 
B7 80 FF FF B3 D1 20 00 13 02 12 00 93 02 20 00 
E3 16 52 FE B7 CE FF 7F 13 0E 20 02 63 9A D1 15 
13 02 00 00 13 01 70 00 B7 80 FF FF 13 00 00 00 
B3 D1 20 00 13 02 12 00 93 02 20 00 E3 14 52 FE 
B7 0E 00 02 93 8E 0E F0 13 0E 30 02 63 92 D1 13 
13 02 00 00 13 01 F0 00 B7 80 FF FF 13 00 00 00 
13 00 00 00 B3 D1 20 00 13 02 12 00 93 02 20 00 
E3 12 52 FE B7 0E 02 00 93 8E FE FF 13 0E 40 02 
63 98 D1 0F 13 02 00 00 13 01 10 00 13 00 00 00 
B7 80 FF FF B3 D1 20 00 13 02 12 00 93 02 20 00 
E3 14 52 FE B7 CE FF 7F 13 0E 50 02 63 92 D1 0D 
13 02 00 00 13 01 70 00 13 00 00 00 B7 80 FF FF 
13 00 00 00 B3 D1 20 00 13 02 12 00 93 02 20 00 
E3 12 52 FE B7 0E 00 02 93 8E 0E F0 13 0E 60 02 
63 98 D1 09 13 02 00 00 13 01 F0 00 13 00 00 00 
13 00 00 00 B7 80 FF FF B3 D1 20 00 13 02 12 00 
93 02 20 00 E3 12 52 FE B7 0E 02 00 93 8E FE FF 
13 0E 70 02 63 9E D1 05 93 00 F0 00 33 51 10 00 
93 0E 00 00 13 0E 80 02 63 14 D1 05 93 00 00 02 
33 D1 00 00 93 0E 00 02 13 0E 90 02 63 1A D1 03 
B3 50 00 00 93 0E 00 00 13 0E A0 02 63 92 D0 03 
93 00 00 40 37 11 00 00 13 01 01 80 33 D0 20 00 
93 0E 00 00 13 0E B0 02 63 14 D0 01 63 1A C0 03 
37 05 00 10 93 05 50 04 13 06 20 05 93 06 F0 04 
13 07 A0 00 23 20 B5 00 23 20 C5 00 23 20 C5 00 
23 20 D5 00 23 20 C5 00 23 20 E5 00 73 00 10 00 
37 05 00 10 93 05 F0 04 13 06 B0 04 93 06 A0 00 
23 20 B5 00 23 20 C5 00 23 20 D5 00 6F F0 5F 9C 
@00000640
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
