`include "rvga_types.svh"

module execute_stage
  ( input logic clk
    , input logic rst
    );

always_ff @(posedge clk) begin

end

always_comb begin

end

endmodule : execute_stage
