@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
