`include "rvga_types.svh"

module decode_stage
(
    input logic clk,
    input logic rst,
    
    input rvga_word ifetch_decode_instruction
);

always_ff @(posedge clk) begin

end

always_comb begin

end

endmodule : decode_stage
