@00000000
37 05 00 00 13 05 05 00 37 06 00 10 83 05 05 00 
63 8C 05 00 23 20 B6 00 13 05 15 00 6F F0 1F FF 
6D 79 74 65 73 74 00 00 93 05 E0 02 23 20 B6 00 
23 20 B6 00 93 00 00 00 13 01 00 00 B3 91 20 02 
93 0E 00 00 13 0E 20 00 63 9A D1 4B 93 00 10 00 
13 01 10 00 B3 91 20 02 93 0E 00 00 13 0E 30 00 
63 9E D1 49 93 00 30 00 13 01 70 00 B3 91 20 02 
93 0E 00 00 13 0E 40 00 63 92 D1 49 93 00 00 00 
37 81 FF FF B3 91 20 02 93 0E 00 00 13 0E 50 00 
63 96 D1 47 B7 00 00 80 13 01 00 00 B3 91 20 02 
93 0E 00 00 13 0E 60 00 63 9A D1 45 B7 00 00 80 
13 01 00 00 B3 91 20 02 93 0E 00 00 13 0E 70 00 
63 9E D1 43 B7 B0 AA AA 93 80 B0 AA 37 01 03 00 
13 01 D1 E7 B3 91 20 02 B7 0E FF FF 93 8E 1E 08 
13 0E E0 01 63 9C D1 41 B7 00 03 00 93 80 D0 E7 
37 B1 AA AA 13 01 B1 AA B3 91 20 02 B7 0E FF FF 
93 8E 1E 08 13 0E F0 01 63 9A D1 3F B7 00 00 FF 
37 01 00 FF B3 91 20 02 B7 0E 01 00 13 0E 00 02 
63 9E D1 3D 93 00 F0 FF 13 01 F0 FF B3 91 20 02 
93 0E 00 00 13 0E 10 02 63 92 D1 3D 93 00 F0 FF 
13 01 10 00 B3 91 20 02 93 0E F0 FF 13 0E 20 02 
63 96 D1 3B 93 00 10 00 13 01 F0 FF B3 91 20 02 
93 0E F0 FF 13 0E 30 02 63 9A D1 39 B7 00 D0 00 
37 01 B0 00 B3 90 20 02 B7 9E 00 00 93 8E 0E F0 
13 0E 80 00 63 9C D0 37 B7 00 E0 00 37 01 B0 00 
33 91 20 02 B7 AE 00 00 93 8E 0E A0 13 0E 90 00 
63 1E D1 35 B7 00 D0 00 B3 90 10 02 B7 BE 00 00 
93 8E 0E 90 13 0E A0 00 63 92 D0 35 13 02 00 00 
B7 00 D0 00 37 01 B0 00 B3 91 20 02 13 83 01 00 
13 02 12 00 93 02 20 00 E3 14 52 FE B7 9E 00 00 
93 8E 0E F0 13 0E B0 00 63 1A D3 31 13 02 00 00 
B7 00 E0 00 37 01 B0 00 B3 91 20 02 13 00 00 00 
13 83 01 00 13 02 12 00 93 02 20 00 E3 12 52 FE 
B7 AE 00 00 93 8E 0E A0 13 0E C0 00 63 10 D3 2F 
13 02 00 00 B7 00 F0 00 37 01 B0 00 B3 91 20 02 
13 00 00 00 13 00 00 00 13 83 01 00 13 02 12 00 
93 02 20 00 E3 10 52 FE B7 AE 00 00 93 8E 0E 50 
13 0E D0 00 63 14 D3 2B 13 02 00 00 B7 00 D0 00 
37 01 B0 00 B3 91 20 02 13 02 12 00 93 02 20 00 
E3 16 52 FE B7 9E 00 00 93 8E 0E F0 13 0E E0 00 
63 9E D1 27 13 02 00 00 B7 00 E0 00 37 01 B0 00 
13 00 00 00 B3 91 20 02 13 02 12 00 93 02 20 00 
E3 14 52 FE B7 AE 00 00 93 8E 0E A0 13 0E F0 00 
63 96 D1 25 13 02 00 00 B7 00 F0 00 37 01 B0 00 
13 00 00 00 13 00 00 00 B3 91 20 02 13 02 12 00 
93 02 20 00 E3 12 52 FE B7 AE 00 00 93 8E 0E 50 
13 0E 00 01 63 9C D1 21 13 02 00 00 B7 00 D0 00 
13 00 00 00 37 01 B0 00 B3 91 20 02 13 02 12 00 
93 02 20 00 E3 14 52 FE B7 9E 00 00 93 8E 0E F0 
13 0E 10 01 63 94 D1 1F 13 02 00 00 B7 00 E0 00 
13 00 00 00 37 01 B0 00 13 00 00 00 B3 91 20 02 
13 02 12 00 93 02 20 00 E3 12 52 FE B7 AE 00 00 
93 8E 0E A0 13 0E 20 01 63 9A D1 1B 13 02 00 00 
B7 00 F0 00 13 00 00 00 13 00 00 00 37 01 B0 00 
B3 91 20 02 13 02 12 00 93 02 20 00 E3 12 52 FE 
B7 AE 00 00 93 8E 0E 50 13 0E 30 01 63 90 D1 19 
13 02 00 00 37 01 B0 00 B7 00 D0 00 B3 91 20 02 
13 02 12 00 93 02 20 00 E3 16 52 FE B7 9E 00 00 
93 8E 0E F0 13 0E 40 01 63 9A D1 15 13 02 00 00 
37 01 B0 00 B7 00 E0 00 13 00 00 00 B3 91 20 02 
13 02 12 00 93 02 20 00 E3 14 52 FE B7 AE 00 00 
93 8E 0E A0 13 0E 50 01 63 92 D1 13 13 02 00 00 
37 01 B0 00 B7 00 F0 00 13 00 00 00 13 00 00 00 
B3 91 20 02 13 02 12 00 93 02 20 00 E3 12 52 FE 
B7 AE 00 00 93 8E 0E 50 13 0E 60 01 63 98 D1 0F 
13 02 00 00 37 01 B0 00 13 00 00 00 B7 00 D0 00 
B3 91 20 02 13 02 12 00 93 02 20 00 E3 14 52 FE 
B7 9E 00 00 93 8E 0E F0 13 0E 70 01 63 90 D1 0D 
13 02 00 00 37 01 B0 00 13 00 00 00 B7 00 E0 00 
13 00 00 00 B3 91 20 02 13 02 12 00 93 02 20 00 
E3 12 52 FE B7 AE 00 00 93 8E 0E A0 13 0E 80 01 
63 96 D1 09 13 02 00 00 37 01 B0 00 13 00 00 00 
13 00 00 00 B7 00 F0 00 B3 91 20 02 13 02 12 00 
93 02 20 00 E3 12 52 FE B7 AE 00 00 93 8E 0E 50 
13 0E 90 01 63 9C D1 05 B7 00 00 7C 33 11 10 02 
93 0E 00 00 13 0E A0 01 63 12 D1 05 B7 00 00 80 
33 91 00 02 93 0E 00 00 13 0E B0 01 63 18 D1 03 
B3 10 00 02 93 0E 00 00 13 0E C0 01 63 90 D0 03 
B7 00 10 02 37 01 20 02 33 90 20 02 93 0E 00 00 
13 0E D0 01 63 14 D0 01 63 1A C0 03 37 05 00 10 
93 05 50 04 13 06 20 05 93 06 F0 04 13 07 A0 00 
23 20 B5 00 23 20 C5 00 23 20 C5 00 23 20 D5 00 
23 20 C5 00 23 20 E5 00 73 00 10 00 37 05 00 10 
93 05 F0 04 13 06 B0 04 93 06 A0 00 23 20 B5 00 
23 20 C5 00 23 20 D5 00 6F F0 9F AB 
@0000054C
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 
