`include "rvga_types.sv"
import rvga_types::*;

`ifndef DEBUG_DEFINES_SVH
`define DEBUG_DEFINES_SVH 1
  `define INST_DEBUG_BUS 1

  `define INST_TRACE_DEBUG 1

  //`define IFETCH_DEBUG
  //`define DECODE_DEBUG
  //`define RFETCH_DEBUG
  //`define EXECUTE_DEBUG
  //`define MEMORY_DEBUG
  //`define WRITEBACK_DEBUG
`endif