@00000000
37 05 00 00 13 05 05 00 37 06 00 10 83 05 05 00 
63 8C 05 00 23 20 B6 00 13 05 15 00 6F F0 1F FF 
6D 79 74 65 73 74 00 00 93 05 E0 02 23 20 B6 00 
23 20 B6 00 97 00 00 00 93 80 00 00 37 01 AA 00 
13 01 A1 0A 23 A0 20 00 83 A1 00 00 B7 0E AA 00 
93 8E AE 0A 13 0E 20 00 63 90 D1 47 97 00 00 00 
93 80 00 00 37 B1 00 AA 13 01 01 A0 23 A2 20 00 
83 A1 40 00 B7 BE 00 AA 93 8E 0E A0 13 0E 30 00 
63 9C D1 43 97 00 00 00 93 80 00 00 37 11 A0 0A 
13 01 01 AA 23 A4 20 00 83 A1 80 00 B7 1E A0 0A 
93 8E 0E AA 13 0E 40 00 63 98 D1 41 97 00 00 00 
93 80 00 00 37 A1 0A A0 13 01 A1 00 23 A6 20 00 
83 A1 C0 00 B7 AE 0A A0 93 8E AE 00 13 0E 50 00 
63 94 D1 3F 97 00 00 00 93 80 00 00 37 01 AA 00 
13 01 A1 0A 23 AA 20 FE 83 A1 40 FF B7 0E AA 00 
93 8E AE 0A 13 0E 60 00 63 90 D1 3D 97 00 00 00 
93 80 00 00 37 B1 00 AA 13 01 01 A0 23 AC 20 FE 
83 A1 80 FF B7 BE 00 AA 93 8E 0E A0 13 0E 70 00 
63 9C D1 39 97 00 00 00 93 80 00 00 37 11 A0 0A 
13 01 01 AA 23 AE 20 FE 83 A1 C0 FF B7 1E A0 0A 
93 8E 0E AA 13 0E 80 00 63 98 D1 37 97 00 00 00 
93 80 00 00 37 A1 0A A0 13 01 A1 00 23 A0 20 00 
83 A1 00 00 B7 AE 0A A0 93 8E AE 00 13 0E 90 00 
63 94 D1 35 97 00 00 00 93 80 00 00 37 51 34 12 
13 01 81 67 13 82 00 FE 23 20 22 02 83 A1 00 00 
B7 5E 34 12 93 8E 8E 67 13 0E A0 00 63 9E D1 31 
97 00 00 00 93 80 00 00 37 31 21 58 13 01 81 09 
93 80 D0 FF A3 A3 20 00 17 02 00 00 13 02 02 00 
83 21 02 00 B7 3E 21 58 93 8E 8E 09 13 0E B0 00 
63 94 D1 2F 13 0E C0 00 13 02 00 00 B7 D0 BB AA 
93 80 D0 CD 17 01 00 00 13 01 01 00 23 20 11 00 
83 21 01 00 B7 DE BB AA 93 8E DE CD 63 9E D1 2B 
13 02 12 00 93 02 20 00 E3 1A 52 FC 13 0E D0 00 
13 02 00 00 B7 C0 AB DA 93 80 D0 CC 17 01 00 00 
13 01 01 00 13 00 00 00 23 22 11 00 83 21 41 00 
B7 CE AB DA 93 8E DE CC 63 90 D1 29 13 02 12 00 
93 02 20 00 E3 18 52 FC 13 0E E0 00 13 02 00 00 
B7 C0 AA DD 93 80 C0 BC 17 01 00 00 13 01 01 00 
13 00 00 00 13 00 00 00 23 24 11 00 83 21 81 00 
B7 CE AA DD 93 8E CE BC 63 90 D1 25 13 02 12 00 
93 02 20 00 E3 16 52 FC 13 0E F0 00 13 02 00 00 
B7 B0 DA CD 93 80 C0 BB 13 00 00 00 17 01 00 00 
13 01 01 00 23 26 11 00 83 21 C1 00 B7 BE DA CD 
93 8E CE BB 63 92 D1 21 13 02 12 00 93 02 20 00 
E3 18 52 FC 13 0E 00 01 13 02 00 00 B7 B0 DD CC 
93 80 B0 AB 13 00 00 00 17 01 00 00 13 01 01 00 
13 00 00 00 23 28 11 00 83 21 01 01 B7 BE DD CC 
93 8E BE AB 63 92 D1 1D 13 02 12 00 93 02 20 00 
E3 16 52 FC 13 0E 10 01 13 02 00 00 B7 E0 CD BC 
93 80 B0 AA 13 00 00 00 13 00 00 00 17 01 00 00 
13 01 01 00 23 2A 11 00 83 21 41 01 B7 EE CD BC 
93 8E BE AA 63 92 D1 19 13 02 12 00 93 02 20 00 
E3 16 52 FC 13 0E 20 01 13 02 00 00 17 01 00 00 
13 01 01 00 B7 20 11 00 93 80 30 23 23 20 11 00 
83 21 01 00 B7 2E 11 00 93 8E 3E 23 63 96 D1 15 
13 02 12 00 93 02 20 00 E3 1A 52 FC 13 0E 30 01 
13 02 00 00 17 01 00 00 13 01 01 00 B7 10 01 30 
93 80 30 22 13 00 00 00 23 22 11 00 83 21 41 00 
B7 1E 01 30 93 8E 3E 22 63 98 D1 11 13 02 12 00 
93 02 20 00 E3 18 52 FC 13 0E 40 01 13 02 00 00 
17 01 00 00 13 01 01 00 B7 10 00 33 93 80 20 12 
13 00 00 00 13 00 00 00 23 24 11 00 83 21 81 00 
B7 1E 00 33 93 8E 2E 12 63 98 D1 0D 13 02 12 00 
93 02 20 00 E3 16 52 FC 13 0E 50 01 13 02 00 00 
17 01 00 00 13 01 01 00 13 00 00 00 B7 00 30 23 
93 80 20 11 23 26 11 00 83 21 C1 00 B7 0E 30 23 
93 8E 2E 11 63 9A D1 09 13 02 12 00 93 02 20 00 
E3 18 52 FC 13 0E 60 01 13 02 00 00 17 01 00 00 
13 01 01 00 13 00 00 00 B7 00 33 22 93 80 10 01 
13 00 00 00 23 28 11 00 83 21 01 01 B7 0E 33 22 
93 8E 1E 01 63 9A D1 05 13 02 12 00 93 02 20 00 
E3 16 52 FC 13 0E 70 01 13 02 00 00 17 01 00 00 
13 01 01 00 13 00 00 00 13 00 00 00 B7 30 23 12 
93 80 10 00 23 2A 11 00 83 21 41 01 B7 3E 23 12 
93 8E 1E 00 63 9A D1 01 13 02 12 00 93 02 20 00 
E3 16 52 FC 63 1A C0 03 37 05 00 10 93 05 50 04 
13 06 20 05 93 06 F0 04 13 07 A0 00 23 20 B5 00 
23 20 C5 00 23 20 C5 00 23 20 D5 00 23 20 C5 00 
23 20 E5 00 73 00 10 00 37 05 00 10 93 05 F0 04 
13 06 B0 04 93 06 A0 00 23 20 B5 00 23 20 C5 00 
23 20 D5 00 6F F0 DF AF 
@00000000
EF BE AD DE EF BE AD DE EF BE AD DE EF BE AD DE 
EF BE AD DE EF BE AD DE EF BE AD DE EF BE AD DE 
EF BE AD DE EF BE AD DE 
@00000508
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 
