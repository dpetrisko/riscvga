@00000000
37 05 00 00 13 05 05 00 37 06 00 10 83 05 05 00 
63 8C 05 00 23 20 B6 00 13 05 15 00 6F F0 1F FF 
6D 79 74 65 73 74 00 00 93 05 E0 02 23 20 B6 00 
23 20 B6 00 B7 00 01 FF 93 80 00 F0 37 11 0F 0F 
13 01 F1 F0 B3 F1 20 00 B7 1E 00 0F 93 8E 0E F0 
13 0E 20 00 63 9C D1 49 B7 10 F0 0F 93 80 00 FF 
37 F1 F0 F0 13 01 01 0F B3 F1 20 00 B7 0E F0 00 
93 8E 0E 0F 13 0E 30 00 63 9A D1 47 B7 00 FF 00 
93 80 F0 0F 37 11 0F 0F 13 01 F1 F0 B3 F1 20 00 
B7 0E 0F 00 93 8E FE 00 13 0E 40 00 63 98 D1 45 
B7 F0 0F F0 93 80 F0 00 37 F1 F0 F0 13 01 01 0F 
B3 F1 20 00 B7 FE 00 F0 13 0E 50 00 63 98 D1 43 
B7 00 01 FF 93 80 00 F0 37 11 0F 0F 13 01 F1 F0 
B3 F0 20 00 B7 1E 00 0F 93 8E 0E F0 13 0E 60 00 
63 96 D0 41 B7 10 F0 0F 93 80 00 FF 37 F1 F0 F0 
13 01 01 0F 33 F1 20 00 B7 0E F0 00 93 8E 0E 0F 
13 0E 70 00 63 14 D1 3F B7 00 01 FF 93 80 00 F0 
B3 F0 10 00 B7 0E 01 FF 93 8E 0E F0 13 0E 80 00 
63 96 D0 3D 13 02 00 00 B7 00 01 FF 93 80 00 F0 
37 11 0F 0F 13 01 F1 F0 B3 F1 20 00 13 83 01 00 
13 02 12 00 93 02 20 00 E3 10 52 FE B7 1E 00 0F 
93 8E 0E F0 13 0E 90 00 63 1A D3 39 13 02 00 00 
B7 10 F0 0F 93 80 00 FF 37 F1 F0 F0 13 01 01 0F 
B3 F1 20 00 13 00 00 00 13 83 01 00 13 02 12 00 
93 02 20 00 E3 1E 52 FC B7 0E F0 00 93 8E 0E 0F 
13 0E A0 00 63 1C D3 35 13 02 00 00 B7 00 FF 00 
93 80 F0 0F 37 11 0F 0F 13 01 F1 F0 B3 F1 20 00 
13 00 00 00 13 00 00 00 13 83 01 00 13 02 12 00 
93 02 20 00 E3 1C 52 FC B7 0E 0F 00 93 8E FE 00 
13 0E B0 00 63 1C D3 31 13 02 00 00 B7 00 01 FF 
93 80 00 F0 37 11 0F 0F 13 01 F1 F0 B3 F1 20 00 
13 02 12 00 93 02 20 00 E3 12 52 FE B7 1E 00 0F 
93 8E 0E F0 13 0E C0 00 63 92 D1 2F 13 02 00 00 
B7 10 F0 0F 93 80 00 FF 37 F1 F0 F0 13 01 01 0F 
13 00 00 00 B3 F1 20 00 13 02 12 00 93 02 20 00 
E3 10 52 FE B7 0E F0 00 93 8E 0E 0F 13 0E D0 00 
63 96 D1 2B 13 02 00 00 B7 00 FF 00 93 80 F0 0F 
37 11 0F 0F 13 01 F1 F0 13 00 00 00 13 00 00 00 
B3 F1 20 00 13 02 12 00 93 02 20 00 E3 1E 52 FC 
B7 0E 0F 00 93 8E FE 00 13 0E E0 00 63 98 D1 27 
13 02 00 00 B7 00 01 FF 93 80 00 F0 13 00 00 00 
37 11 0F 0F 13 01 F1 F0 B3 F1 20 00 13 02 12 00 
93 02 20 00 E3 10 52 FE B7 1E 00 0F 93 8E 0E F0 
13 0E F0 00 63 9C D1 23 13 02 00 00 B7 10 F0 0F 
93 80 00 FF 13 00 00 00 37 F1 F0 F0 13 01 01 0F 
13 00 00 00 B3 F1 20 00 13 02 12 00 93 02 20 00 
E3 1E 52 FC B7 0E F0 00 93 8E 0E 0F 13 0E 00 01 
63 9E D1 1F 13 02 00 00 B7 00 FF 00 93 80 F0 0F 
13 00 00 00 13 00 00 00 37 11 0F 0F 13 01 F1 F0 
B3 F1 20 00 13 02 12 00 93 02 20 00 E3 1E 52 FC 
B7 0E 0F 00 93 8E FE 00 13 0E 10 01 63 90 D1 1D 
13 02 00 00 37 11 0F 0F 13 01 F1 F0 B7 00 01 FF 
93 80 00 F0 B3 F1 20 00 13 02 12 00 93 02 20 00 
E3 12 52 FE B7 1E 00 0F 93 8E 0E F0 13 0E 20 01 
63 96 D1 19 13 02 00 00 37 F1 F0 F0 13 01 01 0F 
B7 10 F0 0F 93 80 00 FF 13 00 00 00 B3 F1 20 00 
13 02 12 00 93 02 20 00 E3 10 52 FE B7 0E F0 00 
93 8E 0E 0F 13 0E 30 01 63 9A D1 15 13 02 00 00 
37 11 0F 0F 13 01 F1 F0 B7 00 FF 00 93 80 F0 0F 
13 00 00 00 13 00 00 00 B3 F1 20 00 13 02 12 00 
93 02 20 00 E3 1E 52 FC B7 0E 0F 00 93 8E FE 00 
13 0E 40 01 63 9C D1 11 13 02 00 00 37 11 0F 0F 
13 01 F1 F0 13 00 00 00 B7 00 01 FF 93 80 00 F0 
B3 F1 20 00 13 02 12 00 93 02 20 00 E3 10 52 FE 
B7 1E 00 0F 93 8E 0E F0 13 0E 50 01 63 90 D1 0F 
13 02 00 00 37 F1 F0 F0 13 01 01 0F 13 00 00 00 
B7 10 F0 0F 93 80 00 FF 13 00 00 00 B3 F1 20 00 
13 02 12 00 93 02 20 00 E3 1E 52 FC B7 0E F0 00 
93 8E 0E 0F 13 0E 60 01 63 92 D1 0B 13 02 00 00 
37 11 0F 0F 13 01 F1 F0 13 00 00 00 13 00 00 00 
B7 00 FF 00 93 80 F0 0F B3 F1 20 00 13 02 12 00 
93 02 20 00 E3 1E 52 FC B7 0E 0F 00 93 8E FE 00 
13 0E 70 01 63 94 D1 07 B7 00 01 FF 93 80 00 F0 
33 71 10 00 93 0E 00 00 13 0E 80 01 63 18 D1 05 
B7 00 FF 00 93 80 F0 0F 33 F1 00 00 93 0E 00 00 
13 0E 90 01 63 1C D1 03 B3 70 00 00 93 0E 00 00 
13 0E A0 01 63 94 D0 03 B7 10 11 11 93 80 10 11 
37 21 22 22 13 01 21 22 33 F0 20 00 93 0E 00 00 
13 0E B0 01 63 14 D0 01 63 1A C0 03 37 05 00 10 
93 05 50 04 13 06 20 05 93 06 F0 04 13 07 A0 00 
23 20 B5 00 23 20 C5 00 23 20 C5 00 23 20 D5 00 
23 20 C5 00 23 20 E5 00 73 00 10 00 37 05 00 10 
93 05 F0 04 13 06 B0 04 93 06 A0 00 23 20 B5 00 
23 20 C5 00 23 20 D5 00 6F F0 9F AC 
@0000053C
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 
