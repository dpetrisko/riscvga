`include "rvga_types.sv"
import rvga_types::*;

module rvga_top #()
(
    input logic clk_i
    , input logic rst_i
    
    /* Instruction cache interface */
    , output rvga_word imem_addr_o
    , input rvga_word imem_data_i
    , input logic imem_resp_v_i
    
    /* Data cache interface */
	, output logic dmem_r_v_o
    , output logic dmem_w_v_o
    , output rvga_word dmem_addr_o
    , input rvga_word dmem_data_i
    , output rvga_word dmem_data_o
    , input logic dmem_resp_v_i
    
    /* Debug Interface */
    , output rvga_writeback_cword debug_word_o
    , output logic debug_word_v_o
);

rvga_word pc;
rvga_word ir;

logic ifetch_stall_v, decode_stall_v, rfetch_stall_v, execute_stall_v, memory_stall_v, writeback_stall_v;
logic ifetch_flush_v, decode_flush_v, rfetch_flush_v, execute_flush_v, memory_flush_v;
logic decode_br_v, rfetch_br_v, execute_br_v, memory_br_v, writeback_br_v;

rvga_decode_cword decode_cword;
rvga_rfetch_cword rfetch_cword;
rvga_execute_cword execute_cword;
rvga_memory_cword memory_cword;
rvga_writeback_cword writeback_cword;

rvga_word writeback_br_tgt;
logic writeback_btaken;

rvga_reg writeback_rd;
rvga_word writeback_rd_data; 
logic writeback_rd_w_v;

  ifetch_stage ifetch(.clk_i(clk_i)
                      ,.rst_i(rst_i)
                      ,.imem_addr_o(imem_addr_o)
                      ,.imem_data_i(imem_data_i)
                      
                      ,.stall_v_i(ifetch_stall_v)
                      ,.flush_v_i(ifetch_flush_v)
                      
                      ,.pc_o(pc)
                      ,.ir_o(ir)
                      
                      ,.br_tgt_i(writeback_br_tgt)
                      ,.btaken_i(writeback_btaken)
                      );
    
  decode_stage decode(.clk_i(clk_i)
                      ,.rst_i(rst_i)
                      
                      ,.stall_v_i(decode_stall_v)
                      ,.flush_v_i(decode_flush_v)
                      
                      ,.pc_i(pc)
                      ,.ir_i(ir)
                      
                      ,.cword_o(decode_cword)
                      
                      ,.br_v_o(decode_br_v)
                      );
    
  rfetch_stage rfetch(.clk_i(clk_i)
                      ,.rst_i(rst_i)
                      
                      ,.stall_v_i(rfetch_stall_v)
                      ,.flush_v_i(rfetch_flush_v)
                      
                      ,.cword_i(decode_cword)
                      ,.cword_o(rfetch_cword)
                      
                      ,.rd_i(writeback_rd)
                      ,.rd_data_i(writeback_rd_data) 
                      ,.rd_w_v_i(writeback_rd_w_v)
                      
                      ,.br_v_o(rfetch_br_v)
                      );
                      
  execute_stage execute(.clk_i(clk_i)
                        ,.rst_i(rst_i)
                        
                        ,.stall_v_i(execute_stall_v)
                        ,.flush_v_i(execute_flush_v)
                        
                        ,.cword_i(rfetch_cword)
                        ,.cword_o(execute_cword)
                        
                        ,.br_v_o(execute_br_v)
                        );
    
  memory_stage memory(.clk_i(clk_i)
                      ,.rst_i(rst_i)
                      
                      ,.stall_v_i(memory_stall_v)
                      ,.flush_v_i(memory_flush_v)
                      
                      ,.cword_i(execute_cword)
                      ,.cword_o(memory_cword)
                      
                      ,.dmem_r_v_o(dmem_r_v_o)
                      ,.dmem_w_v_o(dmem_w_v_o)
                      ,.dmem_addr_o(dmem_addr_o)
                      ,.dmem_data_i(dmem_data_i)
                      ,.dmem_data_o(dmem_data_o)
                      
                      ,.br_v_o(memory_br_v)
                      );
    
  writeback_stage writeback(.clk_i(clk_i)
                            ,.rst_i(rst_i)
                            
                            ,.stall_v_i(writeback_stall_v)
                            
                            ,.cword_i(memory_cword)
                            ,.cword_o(writeback_cword)
                            
                            ,.br_tgt_o(writeback_br_tgt)
                            ,.btaken_o(writeback_btaken)
                            
                            ,.rd_o(writeback_rd)
                            ,.rd_data_o(writeback_rd_data)
                            ,.rd_w_v_o(writeback_rd_w_v)
                            
                            ,.br_v_o(writeback_br_v)
                            );
                            
  hazard hazard(.imem_read_v_i('1)
                ,.imem_resp_v_i(imem_resp_v_i)
                ,.dmem_read_v_i(dmem_r_v_o)
                ,.dmem_resp_v_i(dmem_resp_v_i)
                
                ,.decode_br_v_i(decode_br_v)
                ,.rfetch_br_v_i(rfetch_br_v)
                ,.execute_br_v_i(execute_br_v)
                ,.memory_br_v_i(memory_br_v)
                ,.writeback_br_v_i(writeback_br_v)
                
                ,.ifetch_flush_v_o(ifetch_flush_v)
                ,.decode_flush_v_o(decode_flush_v)
                ,.rfetch_flush_v_o(rfetch_flush_v)
                ,.execute_flush_v_o(execute_flush_v)
                ,.memory_flush_v_o(memory_flush_v)
                
                ,.ifetch_stall_v_o(ifetch_stall_v)
                ,.decode_stall_v_o(decode_stall_v)
                ,.rfetch_stall_v_o(rfetch_stall_v)
                ,.execute_stall_v_o(execute_stall_v)
                ,.memory_stall_v_o(memory_stall_v)
                ,.writeback_stall_v_o(writeback_stall_v)
                ); 

assign debug_word_o = writeback_cword;
assign debug_word_v_o = ~writeback_stall_v;

endmodule : rvga_top
