@00000000
6F 01 00 01 93 00 E0 0D 13 01 D0 0A E7 01 00 00 
93 0F 10 00 E7 01 81 00 13 0F 20 00 
