`ifndef DEBUG_DEFINES_SVH
`define DEBUG_DEFINES_SVH
    `define INST_DEBUG_BUS

    //`define IFETCH_DEBUG
    //`define DECODE_DEBUG
    //`define RFETCH_DEBUG
    //`define EXECUTE_DEBUG
    //`define MEMORY_DEBUG
    //`define WRITEBACK_DEBUG
    
    typedef logic DEBUG_SIGNAL;
`endif