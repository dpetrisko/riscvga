module writeback_dp #()
  ( input logic clk_i
    , input logic rst_i
    );

endmodule : writeback_dp

