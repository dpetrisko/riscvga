`define DDR_DEBUG 1
//`define IMEM_DEBUG 1
`define IF_DEBUG 1
//`define DEC_DEBUG  1
//`define RF_DEBUG   1
//`define EX_DEBUG   1
//`define DMEM_DEBUG 1
//`define WB_DEBUG   1
//`define RF_DEBUG   1
