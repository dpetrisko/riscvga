@00000000
93 00 10 00 13 81 20 00 93 81 30 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
