@00000000
13 00 00 00 13 00 A0 00 93 00 50 00 13 01 F0 FF 
93 01 31 FF 13 A2 60 00 93 A2 40 00 13 B3 31 FF 
93 B3 01 00 13 F4 10 01 93 E4 10 09 13 C5 D4 0B 
93 15 45 00 13 D6 01 01 93 D6 11 40 37 57 34 12 
97 07 00 00 17 A8 00 00 6F 00 00 00 13 00 00 00 
