parameter NUM_REGS = 32,

parameter BYTES_PER_BYTE = 1,
parameter BYTES_PER_SHORT = 2,
parameter BYTES_PER_WORD = 4,

parameter OP_LUI    = 7'b0110111,
parameter OP_AUIPC  = 7'b0010111,
parameter OP_JAL    = 7'b1101111,
parameter OP_JALR   = 7'b1100111,
parameter OP_BR     = 7'b1100011,
parameter OP_LD     = 7'b0000011,
parameter OP_ST     = 7'b0100011,
parameter OP_IMM    = 7'b0010011,
parameter OP_OP     = 7'b0110011,
parameter OP_FENCE  = 7'b0001111,
parameter OP_SYSTEM = 7'b1110011,

parameter NO_OP = 32'b0,

parameter R0  = 5'b00000,
parameter R1  = 5'b00001,
parameter R2  = 5'b00010,
parameter R3  = 5'b00011,
parameter R4  = 5'b00100,
parameter R5  = 5'b00101,
parameter R6  = 5'b00110,
parameter R7  = 5'b00111,
parameter R8  = 5'b01000,
parameter R9  = 5'b01001,
parameter R10 = 5'b01010,
parameter R11 = 5'b01011,
parameter R12 = 5'b01100,
parameter R13 = 5'b01101,
parameter R14 = 5'b01110,
parameter R15 = 5'b01111,
parameter R16 = 5'b10000,
parameter R17 = 5'b10001,
parameter R18 = 5'b10010,
parameter R19 = 5'b10011,
parameter R20 = 5'b10100,
parameter R21 = 5'b10101,
parameter R22 = 5'b10110,
parameter R23 = 5'b10111,
parameter R24 = 5'b11000,
parameter R25 = 5'b11001,
parameter R26 = 5'b11010,
parameter R27 = 5'b11011,
parameter R28 = 5'b11100,
parameter R29 = 5'b11101,
parameter R30 = 5'b11110,
parameter R31 = 5'b11111,

parameter FN3_JALR   = 3'b000,
parameter FN3_BEQ    = 3'b000,
parameter FN3_BNE    = 3'b001,
parameter FN3_BLT    = 3'b100,
parameter FN3_BGE    = 3'b101,
parameter FN3_BLTU   = 3'b110,
parameter FN3_BGEU   = 3'b111,
parameter FN3_LB     = 3'b000,
parameter FN3_LH     = 3'b001,
parameter FN3_LW     = 3'b010,
parameter FN3_LBU    = 3'b100,
parameter FN3_LHU    = 3'b101,
parameter FN3_SB     = 3'b000,
parameter FN3_SH     = 3'b001,
parameter FN3_SW     = 3'b010,
parameter FN3_ADDI   = 3'b000,
parameter FN3_SLTI   = 3'b010,
parameter FN3_SLTIU  = 3'b011,
parameter FN3_XORI   = 3'b100,
parameter FN3_ORI    = 3'b110,
parameter FN3_ANDI   = 3'b111,
parameter FN3_SLLI   = 3'b001,
parameter FN3_SRLI   = 3'b101,
parameter FN3_SRAI   = 3'b101,
parameter FN3_ADD    = 3'b000,
parameter FN3_SUB    = 3'b000,
parameter FN3_SLL    = 3'b001,
parameter FN3_SLT    = 3'b010,
parameter FN3_SLTU   = 3'b011,
parameter FN3_XOR    = 3'b100,
parameter FN3_SRL    = 3'b101,
parameter FN3_SRA    = 3'b101,
parameter FN3_OR     = 3'b110,
parameter FN3_AND    = 3'b111,
parameter FN3_FENCE  = 3'b000,
parameter FN3_FENCEI = 3'b001,
parameter FN3_ECALL  = 3'b000,
parameter FN3_EBREAK = 3'b000,
parameter FN3_CSRRW  = 3'b001,
parameter FN3_CSRRS  = 3'b010,
parameter FN3_CSRRC  = 3'b011,
parameter FN3_CSRRWI = 3'b101,
parameter FN3_CSRRSI = 3'b110,
parameter FN3_CSRRCI = 3'b111,

parameter FN7_SLLI = 7'b0000000,
parameter FN7_SRLI = 7'b0000000,
parameter FN7_SRAI = 7'b0100000,
parameter FN7_ADD  = 7'b0000000,
parameter FN7_SUB  = 7'b0100000

