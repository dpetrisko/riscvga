`include "rvga_types.sv"
import rvga_types::*;

module rfetch_stage
  (input logic clk_i
   , input logic rst_i
   );

endmodule : rfetch_stage

