`ifndef RVGA_DEFINES_SVH
`define RVGA_DEFINES_SVH



`endif
