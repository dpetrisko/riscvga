`include "rvga_types.sv"
import rvga_types::*;

module rfetch_stage
  ( input logic clk
    , input logic rst
    );

always_ff @(posedge clk) begin

end

always_comb begin

end

endmodule : rfetch_stage
