@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
B7 40 23 01 93 80 60 05 17 01 00 00 13 01 01 00 
97 01 00 00 93 81 01 00 17 02 00 00 13 02 02 00 
23 20 11 00 23 90 11 00 23 00 12 00 83 22 01 00 
03 A3 01 00 83 23 02 00 03 14 01 00 83 94 01 00 
03 15 02 00 83 05 01 00 03 86 01 00 83 06 02 00 
6F 00 00 00 13 00 00 00 
@00000000
00 00 00 00 00 00 00 00 00 00 00 00 
