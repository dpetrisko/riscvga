@00000000
37 05 00 00 13 05 05 00 37 06 00 10 83 05 05 00 
63 8C 05 00 23 20 B6 00 13 05 15 00 6F F0 1F FF 
6D 79 74 65 73 74 00 00 93 05 E0 02 23 20 B6 00 
23 20 B6 00 93 00 00 00 13 01 00 00 B3 81 20 40 
93 0E 00 00 13 0E 20 00 63 96 D1 4B 93 00 10 00 
13 01 10 00 B3 81 20 40 93 0E 00 00 13 0E 30 00 
63 9A D1 49 93 00 30 00 13 01 70 00 B3 81 20 40 
93 0E C0 FF 13 0E 40 00 63 9E D1 47 93 00 00 00 
37 81 FF FF B3 81 20 40 B7 8E 00 00 13 0E 50 00 
63 92 D1 47 B7 00 00 80 13 01 00 00 B3 81 20 40 
B7 0E 00 80 13 0E 60 00 63 96 D1 45 B7 00 00 80 
37 81 FF FF B3 81 20 40 B7 8E 00 80 13 0E 70 00 
63 9A D1 43 93 00 00 00 37 81 00 00 13 01 F1 FF 
B3 81 20 40 B7 8E FF FF 93 8E 1E 00 13 0E 80 00 
63 9A D1 41 B7 00 00 80 93 80 F0 FF 13 01 00 00 
B3 81 20 40 B7 0E 00 80 93 8E FE FF 13 0E 90 00 
63 9A D1 3F B7 00 00 80 93 80 F0 FF 37 81 00 00 
13 01 F1 FF B3 81 20 40 B7 8E FF 7F 13 0E A0 00 
63 9A D1 3D B7 00 00 80 37 81 00 00 13 01 F1 FF 
B3 81 20 40 B7 8E FF 7F 93 8E 1E 00 13 0E B0 00 
63 9A D1 3B B7 00 00 80 93 80 F0 FF 37 81 FF FF 
B3 81 20 40 B7 8E 00 80 93 8E FE FF 13 0E C0 00 
63 9A D1 39 93 00 00 00 13 01 F0 FF B3 81 20 40 
93 0E 10 00 13 0E D0 00 63 9E D1 37 93 00 F0 FF 
13 01 10 00 B3 81 20 40 93 0E E0 FF 13 0E E0 00 
63 92 D1 37 93 00 F0 FF 13 01 F0 FF B3 81 20 40 
93 0E 00 00 13 0E F0 00 63 96 D1 35 93 00 D0 00 
13 01 B0 00 B3 80 20 40 93 0E 20 00 13 0E 00 01 
63 9A D0 33 93 00 E0 00 13 01 B0 00 33 81 20 40 
93 0E 30 00 13 0E 10 01 63 1E D1 31 93 00 D0 00 
B3 80 10 40 93 0E 00 00 13 0E 20 01 63 94 D0 31 
13 02 00 00 93 00 D0 00 13 01 B0 00 B3 81 20 40 
13 83 01 00 13 02 12 00 93 02 20 00 E3 14 52 FE 
93 0E 20 00 13 0E 30 01 63 1E D3 2D 13 02 00 00 
93 00 E0 00 13 01 B0 00 B3 81 20 40 13 00 00 00 
13 83 01 00 13 02 12 00 93 02 20 00 E3 12 52 FE 
93 0E 30 00 13 0E 40 01 63 16 D3 2B 13 02 00 00 
93 00 F0 00 13 01 B0 00 B3 81 20 40 13 00 00 00 
13 00 00 00 13 83 01 00 13 02 12 00 93 02 20 00 
E3 10 52 FE 93 0E 40 00 13 0E 50 01 63 1C D3 27 
13 02 00 00 93 00 D0 00 13 01 B0 00 B3 81 20 40 
13 02 12 00 93 02 20 00 E3 16 52 FE 93 0E 20 00 
13 0E 60 01 63 98 D1 25 13 02 00 00 93 00 E0 00 
13 01 B0 00 13 00 00 00 B3 81 20 40 13 02 12 00 
93 02 20 00 E3 14 52 FE 93 0E 30 00 13 0E 70 01 
63 92 D1 23 13 02 00 00 93 00 F0 00 13 01 B0 00 
13 00 00 00 13 00 00 00 B3 81 20 40 13 02 12 00 
93 02 20 00 E3 12 52 FE 93 0E 40 00 13 0E 80 01 
63 9A D1 1F 13 02 00 00 93 00 D0 00 13 00 00 00 
13 01 B0 00 B3 81 20 40 13 02 12 00 93 02 20 00 
E3 14 52 FE 93 0E 20 00 13 0E 90 01 63 94 D1 1D 
13 02 00 00 93 00 E0 00 13 00 00 00 13 01 B0 00 
13 00 00 00 B3 81 20 40 13 02 12 00 93 02 20 00 
E3 12 52 FE 93 0E 30 00 13 0E A0 01 63 9C D1 19 
13 02 00 00 93 00 F0 00 13 00 00 00 13 00 00 00 
13 01 B0 00 B3 81 20 40 13 02 12 00 93 02 20 00 
E3 12 52 FE 93 0E 40 00 13 0E B0 01 63 94 D1 17 
13 02 00 00 13 01 B0 00 93 00 D0 00 B3 81 20 40 
13 02 12 00 93 02 20 00 E3 16 52 FE 93 0E 20 00 
13 0E C0 01 63 90 D1 15 13 02 00 00 13 01 B0 00 
93 00 E0 00 13 00 00 00 B3 81 20 40 13 02 12 00 
93 02 20 00 E3 14 52 FE 93 0E 30 00 13 0E D0 01 
63 9A D1 11 13 02 00 00 13 01 B0 00 93 00 F0 00 
13 00 00 00 13 00 00 00 B3 81 20 40 13 02 12 00 
93 02 20 00 E3 12 52 FE 93 0E 40 00 13 0E E0 01 
63 92 D1 0F 13 02 00 00 13 01 B0 00 13 00 00 00 
93 00 D0 00 B3 81 20 40 13 02 12 00 93 02 20 00 
E3 14 52 FE 93 0E 20 00 13 0E F0 01 63 9C D1 0B 
13 02 00 00 13 01 B0 00 13 00 00 00 93 00 E0 00 
13 00 00 00 B3 81 20 40 13 02 12 00 93 02 20 00 
E3 12 52 FE 93 0E 30 00 13 0E 00 02 63 94 D1 09 
13 02 00 00 13 01 B0 00 13 00 00 00 13 00 00 00 
93 00 F0 00 B3 81 20 40 13 02 12 00 93 02 20 00 
E3 12 52 FE 93 0E 40 00 13 0E 10 02 63 9C D1 05 
93 00 10 FF 33 01 10 40 93 0E F0 00 13 0E 20 02 
63 12 D1 05 93 00 00 02 33 81 00 40 93 0E 00 02 
13 0E 30 02 63 18 D1 03 B3 00 00 40 93 0E 00 00 
13 0E 40 02 63 90 D0 03 93 00 00 01 13 01 E0 01 
33 80 20 40 93 0E 00 00 13 0E 50 02 63 14 D0 01 
63 1A C0 03 37 05 00 10 93 05 50 04 13 06 20 05 
93 06 F0 04 13 07 A0 00 23 20 B5 00 23 20 C5 00 
23 20 C5 00 23 20 D5 00 23 20 C5 00 23 20 E5 00 
73 00 10 00 37 05 00 10 93 05 F0 04 13 06 B0 04 
93 06 A0 00 23 20 B5 00 23 20 C5 00 23 20 D5 00 
6F F0 1F AC 
@00000544
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 
